interface intf(input logic trigger, clk, reset);
  
  //declaring the signals

  logic [7:0] Wb;
  logic mode_a;
   logic mode_b;
  logic delay_out;
  
endinterface
