module delay_timer(input logic trigger, mode_a, mode_b, clk, reset, [7:0]Wb, output reg delay_out);

reg [7:0]timer = 8'b0; //initially timer=0
reg [1:0]mode;
reg timer_start = 1'b0;
reg timer_reset = 1'b0;
reg out=1'b1;
reg [7:0]pulse_width;
logic trigger_2=1'b0;
logic trigger_1=1'b0;
wire trigger_rise, trigger_fall;
reg [7:0]delay;

always_ff@(posedge clk)
begin
assign mode = {mode_a, mode_b};  //programmable mode selection
assign pulse_width = (2*Wb + 1)/2;  //how much delay must be given after the timer starts
end


always_ff@(posedge clk)
begin
trigger_1<= trigger;
trigger_2<= trigger_1;
end

// track of trigger positive & negative transitions
assign trigger_rise = trigger_1 & (~trigger_2); 
assign trigger_fall = trigger_2 & (~trigger_1);

always_comb
begin
case(mode)
	2'b00: begin 		// one-shot mode
		if (trigger_rise==1 && timer<pulse_width) begin
		out<=0;
		timer_start<=1; 
		timer_reset<=0; 
		delay=end
		else	
		if(timer>=pulse_width)begin
		out<=1; 
		timer_reset<=1;
		timer_start<=0; end
		else 
		if(reset)begin
		out<=1;
		timer_reset<=1;
		timer_start<=0; end
end
	2'b01: begin		//delayed operate mode
		if(trigger_rise==1 && timer<pulse_width)begin
		out<=1;
		timer_start<=1;		
		timer_reset<=0;end
		else	
		if(timer>=pulse_width)begin
		out<=0; 
		timer_reset<=1;
		timer_start<=0; end
		else
		if(trigger_fall==1 || trigger==0) begin
		out<=0;
		timer_start<=0;
		timer_reset<=1;end
		else	
		if(reset)begin
		out<=1;
		timer_reset<=1;
		timer_start<=0; end
end
	2'b10: begin			//delayed release mode
		if(reset)begin
		out<=1;
		timer_reset<=1;
		timer_start<=0; end
		else 
		if(trigger==0 && timer<=pulse_width) begin
		out<=0;
		timer_start<=1;
		timer_reset<=0; end
		else
		if(timer>pulse_width)begin
		out<=1;
		timer_start<=0;
		timer_reset<=1;end
		else
		if(trigger_rise==1 || trigger==1) begin
		out<=0;
		timer_start<=0;
		timer_reset<=1;end
end
	2'b11: begin			//dual delay mode
		if(trigger_rise==1 && timer<=pulse_width)begin
		timer_start<=1;
		timer_reset<=0;end
		else
		if(trigger_fall==1 && timer<=pulse_width)begin
		timer_start<=1;
		timer_reset<=0;end
		else
		if(timer>pulse_width)begin
		out<=trigger;
		timer_start<=0;
		timer_reset<=1;end
end
endcase
end

always_ff@(posedge clk) //To start or reset the Timer
begin
	if(timer_start)
	timer <= timer + 1'b1;
	else
	if(timer_reset)
	timer<=0;
end

always_ff@(posedge clk) // Delay output
begin
if(out)
delay_out<=0;
else
delay_out<=1;#10; 
end
endmodule

